module test_design;
    
endmodule