module test_design(
    clk,
    rst_n,
    en,
    wire,
    data
);

endmodule