module SRAMMemory;

endmodule