interface control_if;
    
endinterface